LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY latch1 IS
	PORT( A : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		Resetn, Clock : IN STD_LOGIC;
		Q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
		
END latch1;

ARCHITECTURE Behavior OF latch1 IS
BEGIN 
	PROCESS(Resetn, Clock)
	BEGIN
		IF Resetn = '1' THEN -- If reset is '0' latch doesnt operate
			Q <= "00000000";
		ELSIF Clock'EVENT AND Clock = '1' THEN -- When clock ticks
			Q <= A; -- Set output to the input
		END IF;
	END PROCESS;
END Behavior;